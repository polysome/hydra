typedef Bit#(9) Addr;
typedef Bit#(9) Data;


